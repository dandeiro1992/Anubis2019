`timescale 1ns / 1ps
module Anubis_tb;
   reg [127:0] data_i;
	reg clk,reset;
	reg[1:0] order;
   wire [127:0] data_o; 

Anubis_2 enc(.data_in(data_i),.clk(clk), .reset(reset),.order(order),.data_out(data_o));

initial 
begin
data_i[127:0]=128'h138b408b6E3C231cEDC05b8132dE786e;
reset=1'b1;
order=2'b00;
clk=1'b0;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
reset=1'b0;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
reset=1'b0;
order=2'b01;
data_i[127:0]=128'h8B9cF140834BB85C483AB8FAabefF33C;
#10  clk =  ! clk;
#10  clk =  ! clk;
order=2'b10;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
//0
data_i[127:0]=128'hB7AB13ef9bb0F4Cc61A6caAcfBC00cDA;
reset=1'b1;
order=2'b00;
clk=1'b0;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
reset=1'b0;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
reset=1'b0;
order=2'b01;
data_i[127:0]=128'h7aFC02C32DA7E0865d236Cf1586E1511;
#10  clk =  ! clk;
#10  clk =  ! clk;
order=2'b10;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
//1
data_i[127:0]=128'h09d26d8129ACFf12CD036A45FC2ddc31;
reset=1'b1;
order=2'b00;
clk=1'b0;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
reset=1'b0;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
reset=1'b0;
order=2'b01;
data_i[127:0]=128'h70d4EBCcC01C3E5be7D475679ae61A58;
#10  clk =  ! clk;
#10  clk =  ! clk;
order=2'b10;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
//2
data_i[127:0]=128'h7F6a90Cdd6c9BeE1fB011423cb794fB3;
reset=1'b1;
order=2'b00;
clk=1'b0;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
reset=1'b0;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
reset=1'b0;
order=2'b01;
data_i[127:0]=128'hD971371e3C48AaB7EABD4D4AaBe3f7E8;
#10  clk =  ! clk;
#10  clk =  ! clk;
order=2'b10;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
//3
data_i[127:0]=128'h23d1F777f7ffcCb4FBDA7A6F7FE599CB;
reset=1'b1;
order=2'b00;
clk=1'b0;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
reset=1'b0;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
reset=1'b0;
order=2'b01;
data_i[127:0]=128'hf35D1d604bAA6261E8aa81ad4c7F3aA2;
#10  clk =  ! clk;
#10  clk =  ! clk;
order=2'b10;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
//4
data_i[127:0]=128'hfA6a7922f9bdFC44B3D95F1Cdd7CEE1D;
reset=1'b1;
order=2'b00;
clk=1'b0;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
reset=1'b0;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
reset=1'b0;
order=2'b01;
data_i[127:0]=128'h3a0B6aFa2bdD95065E4BC5cb7CEACcf3;
#10  clk =  ! clk;
#10  clk =  ! clk;
order=2'b10;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
//5
data_i[127:0]=128'hEC8c79598285EADF9136Eca8DDd7EbA7;
reset=1'b1;
order=2'b00;
clk=1'b0;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
reset=1'b0;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
reset=1'b0;
order=2'b01;
data_i[127:0]=128'hCb23E65bABfA9BfDCe94fcB7ab7dEFdB;
#10  clk =  ! clk;
#10  clk =  ! clk;
order=2'b10;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
//6
end

endmodule
