module Inverter(
	input wire [3:0] in_data_1,
	input wire [3:0] in_data_2,
	input wire [3:0] in_data_3,
	input wire [3:0] in_data_4,
	input wire [3:0] in_data_5,

	output wire [3:0] out_data_1,
	output wire [3:0] out_data_2,
	output wire [3:0] out_data_3,
	output wire [3:0] out_data_4,
	output wire [3:0] out_data_5
);

wire [4:0] x;
wire [4:0] y;
wire [4:0] z;
wire [4:0] v;
wire [4:0] o_x;
wire [4:0] o_y;
wire [4:0] o_z;
wire [4:0] o_v;

// change wiring to match the 5-in 5-out paradigm from internal representation.
assign x = {in_data_1[3], in_data_2[3], in_data_3[3], in_data_4[3], in_data_5[3]};
assign y = {in_data_1[2], in_data_2[2], in_data_3[2], in_data_4[2], in_data_5[2]};
assign z = {in_data_1[1], in_data_2[1], in_data_3[1], in_data_4[1], in_data_5[1]};
assign v = {in_data_1[0], in_data_2[0], in_data_3[0], in_data_4[0], in_data_5[0]};

assign out_data_5 ={o_x[0], o_y[0], o_z[0], o_v[0]};
assign out_data_4 ={o_x[1], o_y[1], o_z[1], o_v[1]};
assign out_data_3 ={o_x[2], o_y[2], o_z[2], o_v[2]};
assign out_data_2 ={o_x[3], o_y[3], o_z[3], o_v[3]};
assign out_data_1 ={o_x[4], o_y[4], o_z[4], o_v[4]};

// o_x = XYZ + XV + X + Y shared

assign o_x[0] = ((x[1] ^ x[2] ^ x[3] ^ x[4]) && 
		 (y[1] ^ y[2] ^ y[3] ^ y[4]) && 
		 (z[1] ^ z[2] ^ z[3] ^ z[4])) ^ 
		((x[1] ^ x[2] ^ x[3] ^ x[4]) && 
		 (v[1] ^ v[2] ^ v[3] ^ v[4])) ^ 
		  x[1] ^ y[1];

assign o_x[1] = ((x[0] && (y[2] ^ y[3] ^ y[4]) && (z[2] ^ z[3] ^ z[4])) ^ 
		 (y[0] && (x[2] ^ x[3] ^ x[4]) && (z[2] ^ z[3] ^ z[4])) ^ 
		 (z[0] && (x[2] ^ x[3] ^ x[4]) && (y[2] ^ y[3] ^ y[4])) ^
		 (x[0] && y[0] && (z[2] ^ z[3] ^ z[4])) ^
		 (x[0] && z[0] && (y[2] ^ y[3] ^ y[4])) ^
		 (y[0] && z[0] && (x[2] ^ x[3] ^ x[4])) ^ 
		 (x[0] && y[0] && z[0])) ^ 
		 (x[0] && (v[2] ^ v[3] ^ v[4])) ^
		 (v[0] && (x[2] ^ x[3] ^ x[4])) ^
		 (x[0] && v[0]) ^
		  x[2] ^ y[2];

assign o_x[2] =  (x[0] && y[0] && z[1]) ^ 
		 (x[0] && y[1] && z[0]) ^ 
		 (x[1] && y[0] && z[0]) ^ 
		 (x[0] && y[1] && z[1]) ^ 
		 (x[1] && y[0] && z[1]) ^ 
		 (x[1] && y[1] && z[0]) ^
		 (x[0] && y[1] && z[3]) ^ 
		 (x[1] && y[0] && z[3]) ^ 
		 (x[0] && y[3] && z[1]) ^ 
		 (x[1] && y[3] && z[0]) ^ 
		 (x[3] && y[0] && z[1]) ^ 
		 (x[3] && y[1] && z[0]) ^
	  	 (x[0] && y[1] && z[4]) ^ 
		 (x[1] && y[0] && z[4]) ^ 
		 (x[0] && y[4] && z[1]) ^ 
		 (x[1] && y[4] && z[0]) ^ 
		 (x[4] && y[0] && z[1]) ^ 
		 (x[4] && y[1] && z[0]) ^
		((x[0] && v[1]) ^ (x[1] && v[0])) ^ 
		  x[3] ^ y[3];


assign o_x[3] = (x[0] && y[1] && z[2]) ^ 
		(x[0] && y[2] && z[1]) ^ 
		(x[1] && y[0] && z[2]) ^ 
		(x[1] && y[2] && z[0]) ^ 
		(x[2] && y[0] && z[1]) ^ 
		(x[2] && y[1] && z[0]) ^
		 x[4] ^ y[4];

assign o_x[4] = x[0] ^ y[0];

// o_y = xyz + xyv + yz + xv + y shared

assign o_y[0] = ((x[1] ^ x[2] ^ x[3] ^ x[4]) && 
		 (y[1] ^ y[2] ^ y[3] ^ y[4]) && 
	  	 (v[1] ^ v[2] ^ v[3] ^ v[4])) ^ 
		((x[1] ^ x[2] ^ x[3] ^ x[4]) && 
		 (y[1] ^ y[2] ^ y[3] ^ y[4]) && 
		 (z[1] ^ z[2] ^ z[3] ^ z[4])) ^ 
		((y[1] ^ y[2] ^ y[3] ^ y[4]) && 
		 (z[1] ^ z[2] ^ z[3] ^ z[4])) ^ 
		((x[1] ^ x[2] ^ x[3] ^ x[4]) && 
		 (v[1] ^ v[2] ^ v[3] ^ v[4])) ^ 
		  y[1];

assign o_y[1] = ((x[0] && (y[2] ^ y[3] ^ y[4]) && (v[2] ^ v[3] ^ v[4])) ^
		 (y[0] && (x[2] ^ x[3] ^ x[4]) && (v[2] ^ v[3] ^ v[4])) ^
		 (v[0] && (x[2] ^ x[3] ^ x[4]) && (y[2] ^ y[3] ^ y[4])) ^
		 (x[0] && y[0] && (v[2] ^ v[3] ^ v[4])) ^
		 (x[0] && v[0] && (y[2] ^ y[3] ^ y[4])) ^
		 (y[0] && v[0] && (x[2] ^ x[3] ^ x[4])) ^
		 (x[0] && y[0] && v[0])) ^
		((x[0] && (y[2] ^ y[3] ^ y[4]) && (z[2] ^ z[3] ^ z[4])) ^
		 (y[0] && (x[2] ^ x[3] ^ x[4]) && (z[2] ^ z[3] ^ z[4])) ^
		 (z[0] && (x[2] ^ x[3] ^ x[4]) && (y[2] ^ y[3] ^ y[4])) ^ 
		 (x[0] && y[0] && (z[2] ^ z[3] ^ z[4])) ^
		 (x[0] && z[0] && (y[2] ^ y[3] ^ y[4])) ^ 
		 (y[0] && z[0] && (x[2] ^ x[3] ^ x[4])) ^
		 (x[0] && y[0] && z[0])) ^ 
		 (y[0] && (z[2] ^ z[3] ^ z[4])) ^
		 (z[0] && (y[2] ^ y[3] ^ y[4])) ^ 
		 (y[0] && z[0]) ^
		 (x[0] && (v[2] ^ v[3] ^ v[4])) ^
		 (v[0] && (x[2] ^ x[3] ^ x[4])) ^
		 (x[0] && v[0]) ^ 
		  y[2];

assign o_y[2] = (x[0] && y[0] && v[1]) ^ 
		(x[0] && y[1] && v[0]) ^ 
		(x[1] && y[0] && v[0]) ^ 
		(x[0] && y[1] && v[1]) ^ 
		(x[1] && y[0] && v[1]) ^ 
		(x[1] && y[1] && v[0]) ^
		(x[0] && y[1] && v[3]) ^ 
		(x[1] && y[0] && v[3]) ^ 
		(x[0] && y[3] && v[1]) ^ 
		(x[1] && y[3] && v[0]) ^ 
		(x[3] && y[0] && v[1]) ^ 
		(x[3] && y[1] && v[0]) ^
		(x[0] && y[1] && v[4]) ^ 
		(x[1] && y[0] && v[4]) ^ 
		(x[0] && y[4] && v[1]) ^ 
		(x[1] && y[4] && v[0]) ^ 
		(x[4] && y[0] && v[1]) ^ 
		(x[4] && y[1] && v[0]) ^	
		(x[0] && y[0] && z[1]) ^ 
		(x[0] && y[1] && z[0]) ^ 
		(x[1] && y[0] && z[0]) ^ 
		(x[0] && y[1] && z[1]) ^ 
		(x[1] && y[0] && z[1]) ^ 
		(x[1] && y[1] && z[0]) ^
		(x[0] && y[1] && z[3]) ^ 
		(x[1] && y[0] && z[3]) ^ 
		(x[0] && y[3] && z[1]) ^ 
		(x[1] && y[3] && z[0]) ^ 
		(x[3] && y[0] && z[1]) ^ 
		(x[3] && y[1] && z[0]) ^
		(x[0] && y[1] && z[4]) ^ 
		(x[1] && y[0] && z[4]) ^ 
		(x[0] && y[4] && z[1]) ^ 
		(x[1] && y[4] && z[0]) ^ 
		(x[4] && y[0] && z[1]) ^ 
		(x[4] && y[1] && z[0]) ^
	       ((x[0] && v[1]) ^ (x[1] && v[0])) ^
	       ((y[0] && z[1]) ^ (y[1] && z[0])) ^
		 y[3];

assign o_y[3] = (x[0] && y[1] && v[2]) ^ 
		(x[0] && y[2] && v[1]) ^ 
		(x[1] && y[0] && v[2]) ^ 
		(x[1] && y[2] && v[0]) ^ 
		(x[2] && y[0] && v[1]) ^ 
		(x[2] && y[1] && v[0]) ^
		(x[0] && y[1] && z[2]) ^ 
		(x[0] && y[2] && z[1]) ^ 
		(x[1] && y[0] && z[2]) ^ 
		(x[1] && y[2] && z[0]) ^ 
		(x[2] && y[0] && z[1]) ^ 
		(x[2] && y[1] && z[0]) ^
		 y[4];

assign o_y[4] = y[0];

// XYZ + XZV + YV + Z + Y + X

assign o_z[0] = ((x[1] ^ x[2] ^ x[3] ^ x[4]) && 
		 (y[1] ^ y[2] ^ y[3] ^ y[4]) && 
		 (z[1] ^ z[2] ^ z[3] ^ z[4])) ^ 
		((x[1] ^ x[2] ^ x[3] ^ x[4]) && 
		 (z[1] ^ z[2] ^ z[3] ^ z[4]) && 
		 (v[1] ^ v[2] ^ v[3] ^ v[4])) ^ 
		((y[1] ^ y[2] ^ y[3] ^ y[4]) && 
		 (v[1] ^ v[2] ^ v[3] ^ v[4])) ^ 
		  x[1] ^ y[1] ^ z[1];

assign o_z[1] = ((x[0] && (y[2] ^ y[3] ^ y[4]) && (z[2] ^ z[3] ^ z[4])) ^ 
		 (y[0] && (x[2] ^ x[3] ^ x[4]) && (z[2] ^ z[3] ^ z[4])) ^ 
		 (z[0] && (x[2] ^ x[3] ^ x[4]) && (y[2] ^ y[3] ^ y[4])) ^
		 (x[0] && y[0] && (z[2] ^ z[3] ^ z[4])) ^
		 (x[0] && z[0] && (y[2] ^ y[3] ^ y[4])) ^
		 (y[0] && z[0] && (x[2] ^ x[3] ^ x[4])) ^ 
		 (x[0] && y[0] && z[0])) ^ 
		((x[0] && (z[2] ^ z[3] ^ z[4]) && (v[2] ^ v[3] ^ v[4])) ^ 
		 (z[0] && (x[2] ^ x[3] ^ x[4]) && (v[2] ^ v[3] ^ v[4])) ^ 
		 (v[0] && (x[2] ^ x[3] ^ x[4]) && (z[2] ^ z[3] ^ z[4])) ^
		 (x[0] && z[0] && (v[2] ^ v[3] ^ v[4])) ^
		 (x[0] && v[0] && (z[2] ^ z[3] ^ z[4])) ^
		 (z[0] && v[0] && (x[2] ^ x[3] ^ x[4])) ^ 
		 (x[0] && z[0] && v[0])) ^ 
		 (y[0] && (v[2] ^ v[3] ^ v[4])) ^
		 (v[0] && (y[2] ^ y[3] ^ y[4])) ^
		 (y[0] && v[0]) ^
		  x[2] ^ y[2] ^ z[2];

assign o_z[2] = (x[0] && y[0] && z[1]) ^ 
		(x[0] && y[1] && z[0]) ^ 
		(x[1] && y[0] && z[0]) ^ 
		(x[0] && y[1] && z[1]) ^ 
		(x[1] && y[0] && z[1]) ^ 
		(x[1] && y[1] && z[0]) ^
		(x[0] && y[1] && z[3]) ^ 
		(x[1] && y[0] && z[3]) ^ 
		(x[0] && y[3] && z[1]) ^ 
		(x[1] && y[3] && z[0]) ^ 
		(x[3] && y[0] && z[1]) ^ 
		(x[3] && y[1] && z[0]) ^
		(x[0] && y[1] && z[4]) ^ 
		(x[1] && y[0] && z[4]) ^ 
		(x[0] && y[4] && z[1]) ^ 
		(x[1] && y[4] && z[0]) ^ 
		(x[4] && y[0] && z[1]) ^ 
		(x[4] && y[1] && z[0]) ^
		(x[0] && z[0] && v[1]) ^ 
		(x[0] && z[1] && v[0]) ^ 
		(x[1] && z[0] && v[0]) ^ 
		(x[0] && z[1] && v[1]) ^ 
		(x[1] && z[0] && v[1]) ^ 
		(x[1] && z[1] && v[0]) ^
		(x[0] && z[1] && v[3]) ^ 
		(x[1] && z[0] && v[3]) ^ 
		(x[0] && z[3] && v[1]) ^ 
		(x[1] && z[3] && v[0]) ^ 
		(x[3] && z[0] && v[1]) ^ 
		(x[3] && z[1] && v[0]) ^
		(x[0] && z[1] && v[4]) ^ 
		(x[1] && z[0] && v[4]) ^ 
		(x[0] && z[4] && v[1]) ^ 
		(x[1] && z[4] && v[0]) ^ 
		(x[4] && z[0] && v[1]) ^ 
		(x[4] && z[1] && v[0]) ^
	       ((y[0] && v[1]) ^ (y[1] && v[0])) ^
		 x[3] ^ y[3] ^ z[3];

assign o_z[3] =	(x[0] && y[1] && z[2]) ^ 
		(x[0] && y[2] && z[1]) ^ 
		(x[1] && y[0] && z[2]) ^ 
		(x[1] && y[2] && z[0]) ^ 
		(x[2] && y[0] && z[1]) ^ 
		(x[2] && y[1] && z[0]) ^
		(x[0] && z[1] && v[2]) ^ 
		(x[0] && z[2] && v[1]) ^ 
		(x[1] && z[0] && v[2]) ^ 
		(x[1] && z[2] && v[0]) ^ 
		(x[2] && z[0] && v[1]) ^ 
		(x[2] && z[1] && v[0]) ^
		 x[4] ^ y[4] ^ z[4];

assign o_z[4] = x[0] ^ y[0] ^ z[0];

// XYZ + XYV + XZV + YZV + XZ + XV + YZ + V + Z + Y 

assign o_v[0] = ((x[1] ^ x[2] ^ x[3] ^ x[4]) && 
		 (y[1] ^ y[2] ^ y[3] ^ y[4]) && 
		 (z[1] ^ z[2] ^ z[3] ^ z[4])) ^
		((x[1] ^ x[2] ^ x[3] ^ x[4]) && 
		 (y[1] ^ y[2] ^ y[3] ^ y[4]) && 
	  	 (v[1] ^ v[2] ^ v[3] ^ v[4])) ^ 
		((x[1] ^ x[2] ^ x[3] ^ x[4]) && 
		 (z[1] ^ z[2] ^ z[3] ^ z[4]) && 
		 (v[1] ^ v[2] ^ v[3] ^ v[4])) ^ 
		((y[1] ^ y[2] ^ y[3] ^ y[4]) && 
		 (z[1] ^ z[2] ^ z[3] ^ z[4]) && 
		 (v[1] ^ v[2] ^ v[3] ^ v[4])) ^ 
		((x[1] ^ x[2] ^ x[3] ^ x[4]) && 
		 (z[1] ^ z[2] ^ z[3] ^ z[4])) ^ 		
		((x[1] ^ x[2] ^ x[3] ^ x[4]) && 
		 (v[1] ^ v[2] ^ v[3] ^ v[4])) ^ 
		((y[1] ^ y[2] ^ y[3] ^ y[4]) && 
		 (z[1] ^ z[2] ^ z[3] ^ z[4])) ^ 		
		  y[1] ^ z[1] ^ v[1];

assign o_v[1] = ((x[0] && (y[2] ^ y[3] ^ y[4]) && (z[2] ^ z[3] ^ z[4])) ^ 
		 (y[0] && (x[2] ^ x[3] ^ x[4]) && (z[2] ^ z[3] ^ z[4])) ^ 
		 (z[0] && (x[2] ^ x[3] ^ x[4]) && (y[2] ^ y[3] ^ y[4])) ^
		 (x[0] && y[0] && (z[2] ^ z[3] ^ z[4])) ^
		 (x[0] && z[0] && (y[2] ^ y[3] ^ y[4])) ^
		 (y[0] && z[0] && (x[2] ^ x[3] ^ x[4])) ^ 
		 (x[0] && y[0] && z[0])) ^ 
		((x[0] && (y[2] ^ y[3] ^ y[4]) && (v[2] ^ v[3] ^ v[4])) ^
		 (y[0] && (x[2] ^ x[3] ^ x[4]) && (v[2] ^ v[3] ^ v[4])) ^
		 (v[0] && (x[2] ^ x[3] ^ x[4]) && (y[2] ^ y[3] ^ y[4])) ^
		 (x[0] && y[0] && (v[2] ^ v[3] ^ v[4])) ^
		 (x[0] && v[0] && (y[2] ^ y[3] ^ y[4])) ^
		 (y[0] && v[0] && (x[2] ^ x[3] ^ x[4])) ^
		 (x[0] && y[0] && v[0])) ^
		((x[0] && (z[2] ^ z[3] ^ z[4]) && (v[2] ^ v[3] ^ v[4])) ^ 
		 (z[0] && (x[2] ^ x[3] ^ x[4]) && (v[2] ^ v[3] ^ v[4])) ^ 
		 (v[0] && (x[2] ^ x[3] ^ x[4]) && (z[2] ^ z[3] ^ z[4])) ^
		 (x[0] && z[0] && (v[2] ^ v[3] ^ v[4])) ^
		 (x[0] && v[0] && (z[2] ^ z[3] ^ z[4])) ^
		 (z[0] && v[0] && (x[2] ^ x[3] ^ x[4])) ^ 
		 (x[0] && z[0] && v[0])) ^ 
		((y[0] && (z[2] ^ z[3] ^ z[4]) && (v[2] ^ v[3] ^ v[4])) ^ 
		 (z[0] && (y[2] ^ y[3] ^ y[4]) && (v[2] ^ v[3] ^ v[4])) ^ 
		 (v[0] && (y[2] ^ y[3] ^ y[4]) && (z[2] ^ z[3] ^ z[4])) ^
		 (y[0] && z[0] && (v[2] ^ v[3] ^ v[4])) ^
		 (y[0] && v[0] && (z[2] ^ z[3] ^ z[4])) ^
		 (z[0] && v[0] && (y[2] ^ y[3] ^ y[4])) ^ 
		 (y[0] && z[0] && v[0])) ^
		 (x[0] && (z[2] ^ z[3] ^ z[4])) ^
		 (z[0] && (x[2] ^ x[3] ^ x[4])) ^
		 (x[0] && z[0]) ^ 
		 (x[0] && (v[2] ^ v[3] ^ v[4])) ^
		 (v[0] && (x[2] ^ x[3] ^ x[4])) ^
		 (x[0] && v[0]) ^ 
		 (y[0] && (z[2] ^ z[3] ^ z[4])) ^
		 (z[0] && (y[2] ^ y[3] ^ y[4])) ^ 
		 (y[0] && z[0]) ^
		  y[2] ^ z[2] ^ v[2];

assign o_v[2] = (x[0] && y[0] && z[1]) ^ 
		(x[0] && y[1] && z[0]) ^ 
		(x[1] && y[0] && z[0]) ^ 
		(x[0] && y[1] && z[1]) ^ 
		(x[1] && y[0] && z[1]) ^ 
		(x[1] && y[1] && z[0]) ^
		(x[0] && y[1] && z[3]) ^ 
		(x[1] && y[0] && z[3]) ^ 
		(x[0] && y[3] && z[1]) ^ 
		(x[1] && y[3] && z[0]) ^ 
		(x[3] && y[0] && z[1]) ^ 
		(x[3] && y[1] && z[0]) ^
		(x[0] && y[1] && z[4]) ^ 
		(x[1] && y[0] && z[4]) ^ 
		(x[0] && y[4] && z[1]) ^ 
		(x[1] && y[4] && z[0]) ^ 
		(x[4] && y[0] && z[1]) ^ 
		(x[4] && y[1] && z[0]) ^
		(x[0] && y[0] && v[1]) ^ 
		(x[0] && y[1] && v[0]) ^ 
		(x[1] && y[0] && v[0]) ^ 
		(x[0] && y[1] && v[1]) ^ 
		(x[1] && y[0] && v[1]) ^ 
		(x[1] && y[1] && v[0]) ^
		(x[0] && y[1] && v[3]) ^ 
		(x[1] && y[0] && v[3]) ^ 
		(x[0] && y[3] && v[1]) ^ 
		(x[1] && y[3] && v[0]) ^ 
		(x[3] && y[0] && v[1]) ^ 
		(x[3] && y[1] && v[0]) ^
		(x[0] && y[1] && v[4]) ^ 
		(x[1] && y[0] && v[4]) ^ 
		(x[0] && y[4] && v[1]) ^ 
		(x[1] && y[4] && v[0]) ^ 
		(x[4] && y[0] && v[1]) ^ 
		(x[4] && y[1] && v[0]) ^	
		(x[0] && z[0] && v[1]) ^ 
		(x[0] && z[1] && v[0]) ^ 
		(x[1] && z[0] && v[0]) ^ 
		(x[0] && z[1] && v[1]) ^ 
		(x[1] && z[0] && v[1]) ^ 
		(x[1] && z[1] && v[0]) ^
		(x[0] && z[1] && v[3]) ^ 
		(x[1] && z[0] && v[3]) ^ 
		(x[0] && z[3] && v[1]) ^ 
		(x[1] && z[3] && v[0]) ^ 
		(x[3] && z[0] && v[1]) ^ 
		(x[3] && z[1] && v[0]) ^
		(x[0] && z[1] && v[4]) ^ 
		(x[1] && z[0] && v[4]) ^ 
		(x[0] && z[4] && v[1]) ^ 
		(x[1] && z[4] && v[0]) ^ 
		(x[4] && z[0] && v[1]) ^ 
		(x[4] && z[1] && v[0]) ^
		(y[0] && z[0] && v[1]) ^ 
		(y[0] && z[1] && v[0]) ^ 
		(y[1] && z[0] && v[0]) ^ 
		(y[0] && z[1] && v[1]) ^ 
		(y[1] && z[0] && v[1]) ^ 
		(y[1] && z[1] && v[0]) ^
		(y[0] && z[1] && v[3]) ^ 
		(y[1] && z[0] && v[3]) ^ 
		(y[0] && z[3] && v[1]) ^ 
		(y[1] && z[3] && v[0]) ^ 
		(y[3] && z[0] && v[1]) ^ 
		(y[3] && z[1] && v[0]) ^
		(y[0] && z[1] && v[4]) ^ 
		(y[1] && z[0] && v[4]) ^ 
		(y[0] && z[4] && v[1]) ^ 
		(y[1] && z[4] && v[0]) ^ 
		(y[4] && z[0] && v[1]) ^ 
		(y[4] && z[1] && v[0]) ^
	       ((x[0] && z[1]) ^ (x[1] && z[0])) ^
	       ((x[0] && v[1]) ^ (x[1] && v[0])) ^
	       ((y[0] && z[1]) ^ (y[1] && z[0])) ^
		 y[3] ^ z[3] ^ v[3];

assign o_v[3] = (x[0] && y[1] && z[2]) ^ 
		(x[0] && y[2] && z[1]) ^ 
		(x[1] && y[0] && z[2]) ^ 
		(x[1] && y[2] && z[0]) ^ 
		(x[2] && y[0] && z[1]) ^ 
		(x[2] && y[1] && z[0]) ^
		(x[0] && y[1] && v[2]) ^ 
		(x[0] && y[2] && v[1]) ^ 
		(x[1] && y[0] && v[2]) ^ 
		(x[1] && y[2] && v[0]) ^ 
		(x[2] && y[0] && v[1]) ^ 
		(x[2] && y[1] && v[0]) ^
		(x[0] && z[1] && v[2]) ^ 
		(x[0] && z[2] && v[1]) ^ 
		(x[1] && z[0] && v[2]) ^ 
		(x[1] && z[2] && v[0]) ^ 
		(x[2] && z[0] && v[1]) ^ 
		(x[2] && z[1] && v[0]) ^
		(y[0] && z[1] && v[2]) ^ 
		(y[0] && z[2] && v[1]) ^ 
		(y[1] && z[0] && v[2]) ^ 
		(y[1] && z[2] && v[0]) ^ 
		(y[2] && z[0] && v[1]) ^ 
		(y[2] && z[1] && v[0]) ^
		 y[4] ^ z[4] ^ v[4];

assign o_v[4] = y[0] ^ z[0] ^ v[0];

endmodule

