`timescale 1ns / 1ps
module Anubis_tb;
   reg [127:0] data_i;
	reg clk,reset;
	reg[1:0] order;
   wire [127:0] data_o; 

Anubis_2 enc(.data_in(data_i),.clk(clk), .reset(reset),.order(order),.data_out(data_o));

initial 
begin
data_i[127:0]=128'h80000000000000000000000000000000;
reset=1'b1;
order=2'b00;
clk=1'b0;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
reset=1'b0;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
reset=1'b0;
order = 2'b01;
data_i[127:0]=128'h00000000000000000000000000000000;
#10  clk =  ! clk;
#10  clk =  ! clk;
order = 2'b10;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
data_i[127:0]=128'h01010101010101010101010101010101;
reset=1'b1;
order=2'b00;
clk=1'b0;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
reset=1'b0;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
reset=1'b0;
order = 2'b01;
data_i[127:0]=128'h01010101010101010101010101010101;
#10  clk =  ! clk;
#10  clk =  ! clk;
order = 2'b10;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
data_i[127:0]=128'h00000000000000000000000000000000;
reset=1'b1;
order=2'b00;
clk=1'b0;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
reset=1'b0;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
reset=1'b0;
order = 2'b01;
data_i[127:0]=128'h00000000000000000000000000000000;
#10  clk =  ! clk;
#10  clk =  ! clk;
order = 2'b10;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
end

endmodule
