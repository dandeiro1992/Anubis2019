`timescale 1ns / 1ps
module my_encrypt_tb;
   reg [127:0] data_i;
	reg clk,reset;
	reg [1:0] order;
	reg [127 : 0] random_2;
	reg [127 : 0] random_22;
	reg [127 : 0] random_4;
	reg [127 : 0] random_44;
	reg [127 : 0] random_6;
	reg [19:0] random;
   wire [127:0] data_o; 

Anubis_2 enc(.data_in(data_i),.clk(clk), .reset(reset),.order(order),.data_out(data_o),.random_2(random_2),.random_22(random_22),
					.random_4(random_4),.random_44(random_44),.random_6(random_6),.random(random));


initial 
begin
data_i[127:0]=128'h80000000000000000000000000000000;
random_2=128'h12345000000000000000000000000000;
random_22=128'h00001234500000000000000000000000;
random_4=128'h00000000001234500000000000000000;
random_44=128'h00000000000000123450000000000000;
random_6=128'h00000000000000000000123450000000;
random=20'h12345;
reset=1'b1;
order=2'b00;
clk=1'b0;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
reset=1'b0;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
reset=1'b0;
order = 2'b01;
data_i[127:0]=128'h00000000000000000000000000000000;
#10  clk =  ! clk;
#10  clk =  ! clk;
order = 2'b10;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
data_i[127:0]=128'h01010101010101010101010101010101;
reset=1'b1;
order=2'b00;
clk=1'b0;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
reset=1'b0;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
reset=1'b0;
order = 2'b01;
data_i[127:0]=128'h01010101010101010101010101010101;
#10  clk =  ! clk;
#10  clk =  ! clk;
order = 2'b10;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
#10  clk =  ! clk;
end

endmodule
